module Mem_WB_buff     
    #( parameter    
        WbSize  = 4
    )(
    // input rst, 
    input  clk,enable,

    input  [WbSize-1 :0 ] i_WB,
    input  [31:0] i_MemData ,
    input  [15:0] i_alu,
    input  [2:0 ] i_Rdst, 

    output [2: 0] o_WB,
    output [31:0] o_MemData ,
    output [15:0] o_alu,
    output [ 2:0] o_Rdst 
);
    always @(negedge clk) begin
        // if(rst == 1'b1) begin
        //     o_WB  <=       0;
        //     o_Mem <=       0;
        //     o_alu <=       0;
        //     o_Rdst<=       0;
        // end
        // else 
        if(enable == 1'b1) begin
            o_WB       <=  i_WB;
            o_MemData  <=  i_MemData;
            o_alu      <=  i_alu;
            o_Rdst     <=  i_Rdst;
        end
    end
endmodule
