module CTRL_UNIT(
        clk,
        opcode,
        reset,
        CtrlHaz,
        exceptions,
        interrupts,
        signals
 );

        input clk;
        input [6:0] opcode;
        input reset;
        input CtrlHaz;
        input [3:0]exceptions;
        input [2:0]interrupts;
        output reg [40:0]signals;

	reg isReset;

        always @(*)
        begin: ctrl_unit_op
                if(reset)
		begin
                        signals = 41'b00000000011110001001100111000001111100011;
			isReset = 1;
		end
		else if(isReset)
		begin
			signals = 41'b00000000011111000001100111000001111100011;
			isReset = 0;
		end
                else if(exceptions != 0)
                begin
                        case (exceptions)  
                                4'b0001 :    signals = 41'b00000000011100010001100111000001111100011;
                                4'b0010 :    signals = 41'b00000000011100011001100111000001111100011;
                                4'b0100 :    signals = 41'b00000000011111000001100111000001111100011;
                                4'b1000 :    signals = 41'b00000000011111000001100111000001111100011;
                        endcase
                end
                else if(interrupts != 0)
                begin
                        case (interrupts)  
                                3'b001 :    signals = 41'b00000000000000100001100111000001111100011;
                                3'b010 :    signals = 41'b00000000000000101001100111000001111100011;
                                3'b100 :    signals = 41'b00000000011101000001100111000001111100011;
                        endcase
                end
                else
                        case (opcode)  
                                7'b0000000 :    signals = 41'b00000000000000000001100111000001110100001;
                                //one operand
                                7'b0010001 :    signals = 41'b00000000000000000001110111000001001100011; //NOT
                                7'b0000011 :    signals = 41'b00000000000000000001110110000000001100011; //INC
                                7'b0011001 :    signals = 41'b00000000000000000101100111000001011100011; //OUT
                                7'b0011000 :    signals = 41'b00000000000000000001111111000001011100011; //IN
                                7'b1100001 :    signals = 41'b00000000000000000000100111000001111100011; //HLT
                                7'b1101000 :    signals = 41'b00000000000000000001100111000001111100001; //NOP
                                7'b1100010 :    signals = 41'b00000000000000000001100111000000011100011; //SET C
                                //two operand
                                7'b0010101 :    signals = 41'b00000000000000000001110111000001011100011; //MOV
                                7'b0000001 :    signals = 41'b00000000000000000001110111000000001100011; //ADD
                                7'b0001001 :    signals = 41'b00000000000000000001110111000000101100011; //SUB
                                7'b0001101 :    signals = 41'b00000000000000000001110111000000111100011; //AND
                                7'b0100000 :    signals = 41'b00000000000000000010110111100000001100011; //IADD
                                //memory operations
                                7'b0110101 :    signals = 41'b00000000000000000010110111100001101100011; //LDM
                                7'b0100010 :    signals = 41'b00000000000000000010110111100000001110010; //LDD
                                7'b0100011 :    signals = 41'b00000000000000000010100101100000001101011; //STD
                                7'b1110010 :    signals = 41'b00001110000000000001100111000001011101011; //PUSH
                                7'b1110101 :    signals = 41'b00001001100000000001110111000001011110010; //POP
                                //branch operations
                                7'b1010100 :    signals = 41'b00010000000000000001100111000001011100011; //JZ
                                7'b1010101 :    signals = 41'b00100000000000000001100111000001011100011; //JN
                                7'b1010110 :    signals = 41'b00110000000000000001100111000001011100011; //JC
                                7'b1010111 :    signals = 41'b01000000000000000001100111000001011100011; //JMP
                                7'b1111010 :    signals = 41'b11001101000000000001100111000001011101111; //CALL
                                7'b1111110 :    signals = 41'b11001101000000000001100111000001011101111; //INT
                        endcase
                
                if(CtrlHaz)
                begin
                  signals[27:24] = 4'b0111;
                  signals[31:28] = 4'b0100;
                end
        end // ctrl_unit_op
endmodule // CTRL_UNIT